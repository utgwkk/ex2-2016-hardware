* kadai2-1
.include logic.cir
.options post temp=27

v1 in 0 pwl ( 0.0n 0.0
+             4.9n 0.0
+             5.0n 2.5
+             9.9n 2.5
+            10.0n 0.0
+            14.9n 0.0
+            15.0n 2.5)
vdd 1 0 2.5
x1 in out 1 inv
c1 out 0 30f

.tran 0.0005n 20n
.end

* down: 5.013750e-09 - 4.900000e-09 = 1.1375e-10
* up: 1.003025e-08 - 9.900000e-09 = 1.3025e-10
